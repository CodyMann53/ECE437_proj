/*
  Cody Mann
  mann53@purdue.edu

  register file 
*/
